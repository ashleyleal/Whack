// Top Level Module (Main)

module top_module {

}
endmodule